// File: common_defines.svh
`ifndef COMMON_DEFINES_SVH
`define COMMON_DEFINES_SVH

typedef enum {
  CREDIT,
  START,
  EATING_PACDOT,
  EATING_GHOST,
  BLUE_GHOST_MODE,
  GAME_PLAY,
  FAIL,
  FINISH
} sound_t;

`endif
