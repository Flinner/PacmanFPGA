module top_square #(
    parameter CORDW = 10
) (  // coordinate width
    input  wire logic             clk_pix,  // pixel clock
    input  wire logic             sim_rst,  // sim reset
    output logic      [CORDW-1:0] sdl_sx,   // horizontal SDL position
    output logic      [CORDW-1:0] sdl_sy,   // vertical SDL position
    output logic                  sdl_de,   // data enable (low in blanking interval)
    output logic      [      7:0] sdl_r,    // 8-bit red
    output logic      [      7:0] sdl_g,    // 8-bit green
    output logic      [      7:0] sdl_b     // 8-bit blue
);

  // display sync signals and coordinates
  logic [CORDW-1:0] sx, sy;
  logic de;
  simple_480p display_inst (
      .clk_pix,
      .rst_pix(sim_rst),
      .sx,
      .sy,
      .hsync  (),
      .vsync  (),
      .de
  );

  // define a square with screen coordinates
  logic square;
  always_comb begin
    square = (sx > 220 && sx < 420) && (sy > 140 && sy < 340);
  end

  // paint colours: white inside square, blue outside
  logic [3:0] paint_r, paint_g, paint_b;
  always_comb begin
    paint_r = (square) ? 4'hF : 4'h1;
    paint_g = (square) ? 4'hF : 4'h3;
    paint_b = (square) ? 4'hF : 4'h7;
  end

  // SDL output (8 bits per colour channel)
  always_ff @(posedge clk_pix) begin
    sdl_sx <= sx;
    sdl_sy <= sy;
    sdl_de <= de;
    sdl_r  <= {2{paint_r}};  // double signal width from 4 to 8 bits
    sdl_g  <= {2{paint_g}};
    sdl_b  <= {2{paint_b}};
  end
endmodule
